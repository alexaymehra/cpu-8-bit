`timescale 1ns / 1ps
module tb_control_unit_execute;

    reg [7:0] instr;
    reg [2:0] state;
    reg zf;
    reg reset;

    wire [2:0] next_state;
    wire pc_we;
    wire pc_sel;
    wire pc_jmp_sel;
    wire [3:0] pc_offset;
    wire addr_sel;
    wire [3:0] addr_offset;
    wire mem_sel;
    wire mem_we;
    wire [2:0] alu_opcode;
    wire alu_sel_a;
    wire alu_sel_b;
    wire alu_we;
    wire zf_we;
    wire ir_we;
    wire a_sel;
    wire b_sel;
    wire b_we;
    wire halt;

    // FSM States --------------------------------
    localparam FETCH      = 3'b000; 
    localparam DECODE     = 3'b001;
    localparam EXECUTE    = 3'b010;
    localparam MEMORY     = 3'b011;
    localparam WRITEBACK  = 3'b100;
    localparam HALT_STATE = 3'b101;
    localparam IDLE       = 3'b110;
    // -------------------------------------------

    control_unit control_unit_8b (
        .instr(instr),
        .state(state),
        .zf(zf),
        .reset(reset),
        .next_state(next_state),
        .pc_we(pc_we),
        .pc_sel(pc_sel),
        .pc_jmp_sel(pc_jmp_sel),
        .pc_offset(pc_offset),
        .addr_sel(addr_sel),
        .addr_offset(addr_offset),
        .mem_sel(mem_sel),
        .mem_we(mem_we),
        .alu_opcode(alu_opcode),
        .alu_sel_a(alu_sel_a),
        .alu_sel_b(alu_sel_b),
        .alu_we(alu_we),
        .zf_we(zf_we),
        .ir_we(ir_we),
        .a_sel(a_sel),
        .a_we(a_we),
        .b_sel(b_sel),
        .b_we(b_we),
        .halt(halt)
    );

    initial begin
        $dumpfile("control_unitTB_execute.vcd");
        $dumpvars(0, tb_control_unit_execute);
    end

    integer pass_count = 0;
    integer fail_count = 0;

    task automatic check_execute; 
        input integer test_num;
        input [2:0] exp_next_state;
        input [2:0] exp_alu_opcode;
        input exp_alu_sel_a;
        input exp_alu_sel_b;
        input exp_alu_we;
        input exp_zf_we;
        input [3:0] exp_pc_offset;
        input exp_pc_jmp_sel;
        input exp_pc_sel;
        input exp_pc_we;
        integer failed;
    begin
        $display("----- Beginning Test %0d -----", test_num);

        failed = 0;

        if (next_state != exp_next_state) begin
            $display("Test %0d Failed: next_state", test_num);
            failed = 1;
        end

        if (pc_we != exp_pc_we) begin
            $display("Test %0d Failed: pc_we", test_num);
            failed = 1;
        end

        if (pc_sel != exp_pc_sel) begin
            $display("Test %0d Failed: pc_sel", test_num);
            failed = 1;
        end

        if (pc_jmp_sel != exp_pc_jmp_sel) begin
            $display("Test %0d Failed: pc_jmp_sel", test_num);
            failed = 1;
        end

        if (pc_offset != exp_pc_offset) begin
            $display("Test %0d Failed: pc_offset", test_num);
            failed = 1;
        end

        if (addr_sel != 0) begin
            $display("Test %0d Failed: addr_sel", test_num);
            failed = 1;
        end

        if (addr_offset != 4'b0000) begin
            $display("Test %0d Failed: addr_offset", test_num);
            failed = 1;
        end

        if (mem_sel != 0) begin
            $display("Test %0d Failed: mem_sel", test_num);
            failed = 1;
        end

        if (mem_we != 0) begin
            $display("Test %0d Failed: mem_we", test_num);
            failed = 1;
        end

        if (alu_opcode != exp_alu_opcode) begin
            $display("Test %0d Failed: alu_opcode", test_num);
            failed = 1;
        end

        if (alu_sel_a != exp_alu_sel_a) begin
            $display("Test %0d Failed: alu_sel_a", test_num);
            failed = 1;
        end

        if (alu_sel_b != exp_alu_sel_b) begin
            $display("Test %0d Failed: alu_sel_b", test_num);
            failed = 1;
        end

        if (alu_we != exp_alu_we) begin
            $display("Test %0d Failed: alu_we", test_num);
            failed = 1;
        end

        if (zf_we != exp_zf_we) begin
            $display("Test %0d Failed: zf_we", test_num);
            failed = 1;
        end

        if (ir_we != 0) begin
            $display("Test %0d Failed: ir_we", test_num);
            failed = 1;
        end

        if (a_sel != 0) begin
            $display("Test %0d Failed: a_sel", test_num);
            failed = 1;
        end

        if (a_we != 0) begin
            $display("Test %0d Failed: a_we", test_num);
            failed = 1;
        end

        if (b_sel != 0) begin
            $display("Test %0d Failed: b_sel", test_num);
            failed = 1;
        end

        if (b_we != 0) begin
            $display("Test %0d Failed: b_we", test_num);
            failed = 1;
        end

        if (halt != 0) begin
            $display("Test %0d Failed: halt", test_num);
            failed = 1;
        end

        if (failed) begin
            fail_count = fail_count + 1;
            $display("Test %0d RESULT: FAIL\n", test_num);
        end else begin
            pass_count = pass_count + 1;
            $display("Test %0d RESULT: PASS\n", test_num);
        end
    end
    endtask



    initial begin

        // Testing EXECUTE
        $display("Testing EXECUTE\n");
        reset = 1; #10;
        reset = 0; state = EXECUTE; zf = 0;

        instr = 8'b00010100; #10;   // ADD B, A, B
        check_execute(
            1,          // test_num
            WRITEBACK,  // exp_next_state
            3'b000,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b1,       // exp_alu_sel_b
            1'b1,       // exp_alu_we
            1'b1,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        instr = 8'b00001000; #10;   // ADD A, B, A
        check_execute(
            2,          // test_num
            WRITEBACK,  // exp_next_state
            3'b000,     // exp_alu_opcode
            1'b1,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b1,       // exp_alu_we
            1'b1,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        instr = 8'b00110100; #10;   // AND B, A, B
        check_execute(
            3,          // test_num
            WRITEBACK,  // exp_next_state
            3'b001,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b1,       // exp_alu_sel_b
            1'b1,       // exp_alu_we
            1'b1,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        instr = 8'b00101000; #10;   // AND A, B, A
        check_execute(
            4,          // test_num
            WRITEBACK,  // exp_next_state
            3'b001,     // exp_alu_opcode
            1'b1,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b1,       // exp_alu_we
            1'b1,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        instr = 8'b01001000; #10;   // NOT A, B
        check_execute(
            5,          // test_num
            WRITEBACK,  // exp_next_state
            3'b010,     // exp_alu_opcode
            1'b1,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b1,       // exp_alu_we
            1'b1,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        instr = 8'b01010000; #10;   // NOT B, A
        check_execute(
            6,          // test_num
            WRITEBACK,  // exp_next_state
            3'b010,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b1,       // exp_alu_we
            1'b1,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        instr = 8'b10101111; #10;   // JUMP A, 15
        check_execute(
            7,          // test_num
            FETCH,      // exp_next_state
            3'b000,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b0,       // exp_alu_we
            1'b0,       // exp_zf_we
            4'b1111,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b1,       // exp_pc_sel
            1'b1        // exp_pc_we
        );

        instr = 8'b10110101; #10;   // JUMP B, 5
        check_execute(
            8,          // test_num
            FETCH,      // exp_next_state
            3'b000,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b0,       // exp_alu_we
            1'b0,       // exp_zf_we
            4'b0101,    // exp_pc_offset
            1'b1,       // exp_pc_jmp_sel
            1'b1,       // exp_pc_sel
            1'b1        // exp_pc_we
        );

        instr = 8'b11010011; #10;   // JUMPz B, 3 (zf = 0)
        check_execute(
            9,          // test_num
            FETCH,      // exp_next_state
            3'b000,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b0,       // exp_alu_we
            1'b0,       // exp_zf_we
            4'b0000,    // exp_pc_offset
            1'b0,       // exp_pc_jmp_sel
            1'b0,       // exp_pc_sel
            1'b0        // exp_pc_we
        );

        zf = 1; #10;                // JUMPz B, 3 (zf = 1)
        check_execute(
            10,         // test_num
            FETCH,      // exp_next_state
            3'b000,     // exp_alu_opcode
            1'b0,       // exp_alu_sel_a
            1'b0,       // exp_alu_sel_b
            1'b0,       // exp_alu_we
            1'b0,       // exp_zf_we
            4'b0011,    // exp_pc_offset
            1'b1,       // exp_pc_jmp_sel
            1'b1,       // exp_pc_sel
            1'b1        // exp_pc_we
        );

        
        $display("=================================");
        $display("TEST SUMMARY");
        $display("Passed: %0d", pass_count);
        $display("Failed: %0d", fail_count);
        $display("=================================");
        $finish;

    end

endmodule;